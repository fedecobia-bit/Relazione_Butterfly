-- Federico Cobianchi - 332753
-- Onice Mazzi - 359754
-- Antonio Telmon - 353781

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.fixed_float_types.all;
use IEEE.fixed_pkg.all;

entity tb_fft is
end	tb_fft;

architecture behavioral of tb_fft is
	
component BFLY_TOP_ENTITY is
	port(	
		-- segnali reali ingresso
		x0r_in, x1r_in, x2r_in, x3r_in, x4r_in, x5r_in, x6r_in, x7r_in:	in	STD_LOGIC_VECTOR (23 downto 0);
		x8r_in, x9r_in, x10r_in, x11r_in, x12r_in, x13r_in, x14r_in, x15r_in:	in	STD_LOGIC_VECTOR (23 downto 0);
		-- segnali immaginari ingresso
		x0i_in, x1i_in, x2i_in, x3i_in, x4i_in, x5i_in, x6i_in, x7i_in:	in	STD_LOGIC_VECTOR (23 downto 0);
		x8i_in, x9i_in, x10i_in, x11i_in, x12i_in, x13i_in, x14i_in, x15i_in:	in	STD_LOGIC_VECTOR (23 downto 0);
		-- segnali reali uscita
		x0r_out, x1r_out, x2r_out, x3r_out, x4r_out, x5r_out, x6r_out, x7r_out:	out	STD_LOGIC_VECTOR (23 downto 0);
		x8r_out, x9r_out, x10r_out, x11r_out, x12r_out, x13r_out, x14r_out, x15r_out:	out	STD_LOGIC_VECTOR (23 downto 0);
		-- segnali immaginari uscita
		x0i_out, x1i_out, x2i_out, x3i_out, x4i_out, x5i_out, x6i_out, x7i_out:	out	STD_LOGIC_VECTOR (23 downto 0);
		x8i_out, x9i_out, x10i_out, x11i_out, x12i_out, x13i_out, x14i_out, x15i_out:	out	STD_LOGIC_VECTOR (23 downto 0);
		-- segnali di controllo
		Clock: in STD_LOGIC;
		START : in STD_LOGIC;
		DONE : out STD_LOGIC
		);
end component;

	constant period : time := 10 ns; --  clock da 100MHz
	
	signal TB_CLK: STD_LOGIC := '0';
	signal TB_START: STD_LOGIC := '0';
	signal TB_DONE: STD_LOGIC := '0';
	type array_dati is array (0 to 15) of STD_LOGIC_VECTOR(23 downto 0);
   signal r_in : array_dati := (others => (others => '0')); -- other piu' annidato mette tutto a 0, l'altro lo fa per tutte le posizioni
   signal i_in : array_dati := (others => (others => '0'));
   signal r_out : array_dati;
   signal i_out : array_dati;
   
   type sfixed_array is array (0 to 15) of sfixed (0 downto -23);
   
   signal sfixed_xr_in, sfixed_xi_in : sfixed_array;
   signal sfixed_xr_out, sfixed_xi_out : sfixed_array;
   
	
	begin
	
	for_sfixed : for j in 0 to 15 generate
			sfixed_xr_in(j) <= to_sfixed((r_in(j)),0,-23); 
			sfixed_xi_in(j) <= to_sfixed((i_in(j)),0,-23);

			sfixed_xr_out(j) <= to_sfixed((r_out(j)),0,-23);
			sfixed_xi_out(j) <= to_sfixed((i_out(j)),0,-23);

	end generate;
	
	TB_CLK <= not TB_CLK after period/2;
	
	DUT : BFLY_TOP_ENTITY port map (
	-- assegnazione dei segnali di controllo
		Clock => TB_CLK,
		START => TB_START,
		DONE  => TB_DONE,
	-- assegnazione dei segnali ingresso reali
		x0r_in => r_in(0),
		x1r_in => r_in(1),
		x2r_in => r_in(2),
		x3r_in => r_in(3),
		x4r_in => r_in(4),
		x5r_in => r_in(5),
		x6r_in => r_in(6),
		x7r_in => r_in(7),
		x8r_in => r_in(8),
		x9r_in => r_in(9),
		x10r_in => r_in(10),
		x11r_in => r_in(11),
		x12r_in => r_in(12),
		x13r_in => r_in(13),
		x14r_in => r_in(14),
		x15r_in => r_in(15),
	-- assegnazione dei segnali ingresso immaginari
		x0i_in => i_in(0),
		x1i_in => i_in(1),
		x2i_in => i_in(2),
		x3i_in => i_in(3),
		x4i_in => i_in(4),
		x5i_in => i_in(5),
		x6i_in => i_in(6),
		x7i_in => i_in(7),
		x8i_in => i_in(8),
		x9i_in => i_in(9),
		x10i_in => i_in(10),
		x11i_in => i_in(11),
		x12i_in => i_in(12),
		x13i_in => i_in(13),
		x14i_in => i_in(14),
		x15i_in => i_in(15),
	-- assegnazione dei segnali d'uscita reali
		x0r_out => r_out(0),
		x1r_out => r_out(1),
		x2r_out => r_out(2),
		x3r_out => r_out(3),
		x4r_out => r_out(4),
		x5r_out => r_out(5),
		x6r_out => r_out(6),
		x7r_out => r_out(7),
		x8r_out => r_out(8),
		x9r_out => r_out(9),
		x10r_out => r_out(10),
		x11r_out => r_out(11),
		x12r_out => r_out(12),
		x13r_out => r_out(13),
		x14r_out => r_out(14),
		x15r_out => r_out(15),
	-- assegnazione dei segnali d'uscita immaginari
		x0i_out => i_out(0),
		x1i_out => i_out(1),
		x2i_out => i_out(2),
		x3i_out => i_out(3),
		x4i_out => i_out(4),
		x5i_out => i_out(5),
		x6i_out => i_out(6),
		x7i_out => i_out(7),
		x8i_out => i_out(8),
		x9i_out => i_out(9),
		x10i_out => i_out(10),
		x11i_out => i_out(11),
		x12i_out => i_out(12),
		x13i_out => i_out(13),
		x14i_out => i_out(14),
		x15i_out => i_out(15)
    );
	 
	 
	 
	process
    begin
	 TB_START <= '0';
    wait for 2*period; -- Aspetto 2 period prima di iniziare la simulazione
	TB_START <= '1';
	 
	 ---------------------- TEST 1 ----------------------	-1 -1 -1 -1 -1 -1 -1 -1 -1 -1 -1 -1 -1 -1 -1 -1
		r_in(0) <= "100000000000000000000000";
		r_in(1) <= "100000000000000000000000";
		r_in(2) <= "100000000000000000000000";
		r_in(3) <= "100000000000000000000000";
		r_in(4) <= "100000000000000000000000";
		r_in(5) <= "100000000000000000000000";
		r_in(6) <= "100000000000000000000000";
		r_in(7) <= "100000000000000000000000";
		r_in(8) <= "100000000000000000000000";
		r_in(9) <= "100000000000000000000000";
		r_in(10) <= "100000000000000000000000";
		r_in(11) <= "100000000000000000000000";
		r_in(12) <= "100000000000000000000000";
		r_in(13) <= "100000000000000000000000";
		r_in(14) <= "100000000000000000000000";
		r_in(15) <= "100000000000000000000000";
		
		i_in(0) <= "000000000000000000000000";
		i_in(1) <= "000000000000000000000000";
		i_in(2) <= "000000000000000000000000";
		i_in(3) <= "000000000000000000000000";
		i_in(4) <= "000000000000000000000000";
		i_in(5) <= "000000000000000000000000";
		i_in(6) <= "000000000000000000000000";
		i_in(7) <= "000000000000000000000000";
		i_in(8) <= "000000000000000000000000";
		i_in(9) <= "000000000000000000000000";
		i_in(10) <= "000000000000000000000000";
		i_in(11) <= "000000000000000000000000";
		i_in(12) <= "000000000000000000000000";
		i_in(13) <= "000000000000000000000000";
		i_in(14) <= "000000000000000000000000";
		i_in(15) <= "000000000000000000000000";
	 
    wait for 2*period;
    TB_START <= '0';
	
	wait for 11*period;
	TB_START <= '1';
			
	---------------------- TEST 2 ---------------------- -1 0 1 0 -1 0 1 0 -1 0 1 0 -1 0 1 0	
		r_in(0) <= "100000000000000000000000";
		r_in(1) <= "000000000000000000000000";
		r_in(2) <= "011111111111111111111111";
		r_in(3) <= "000000000000000000000000";
		r_in(4) <= "100000000000000000000000";
		r_in(5) <= "000000000000000000000000";
		r_in(6) <= "011111111111111111111111";
		r_in(7) <= "000000000000000000000000";
		r_in(8) <= "100000000000000000000000";
		r_in(9) <= "000000000000000000000000";
		r_in(10) <= "011111111111111111111111";
		r_in(11) <= "000000000000000000000000";
		r_in(12) <= "100000000000000000000000";
		r_in(13) <= "000000000000000000000000";
		r_in(14) <= "011111111111111111111111";
		r_in(15) <= "000000000000000000000000";
		
		i_in(0) <= "000000000000000000000000";
		i_in(1) <= "000000000000000000000000";
		i_in(2) <= "000000000000000000000000";
		i_in(3) <= "000000000000000000000000";
		i_in(4) <= "000000000000000000000000";
		i_in(5) <= "000000000000000000000000";
		i_in(6) <= "000000000000000000000000";
		i_in(7) <= "000000000000000000000000";
		i_in(8) <= "000000000000000000000000";
		i_in(9) <= "000000000000000000000000";
		i_in(10) <= "000000000000000000000000";
		i_in(11) <= "000000000000000000000000";
		i_in(12) <= "000000000000000000000000";
		i_in(13) <= "000000000000000000000000";
		i_in(14) <= "000000000000000000000000";
		i_in(15) <= "000000000000000000000000";
	 
	 wait for 1*period;
	 TB_START <= '0';

	wait for 12*period;
	TB_START <= '1';
			
		---------------------- TEST 3 ----------------------	1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
		 r_in(0) <= "011111111111111111111111";
		 r_in(1) <= "000000000000000000000000";
		 r_in(2) <= "000000000000000000000000";
		 r_in(3) <= "000000000000000000000000";
		 r_in(4) <= "000000000000000000000000";
		 r_in(5) <= "000000000000000000000000";
		 r_in(6) <= "000000000000000000000000";
		 r_in(7) <= "000000000000000000000000";
		 r_in(8) <= "000000000000000000000000";
		 r_in(9) <= "000000000000000000000000";
		 r_in(10) <= "000000000000000000000000";
		 r_in(11) <= "000000000000000000000000";
		 r_in(12) <= "000000000000000000000000";
		 r_in(13) <= "000000000000000000000000";
		 r_in(14) <= "000000000000000000000000";
		 r_in(15) <= "000000000000000000000000";
		 
		 i_in(0) <= "000000000000000000000000";
		 i_in(1) <= "000000000000000000000000";
		 i_in(2) <= "000000000000000000000000";
		 i_in(3) <= "000000000000000000000000";
		 i_in(4) <= "000000000000000000000000";
		 i_in(5) <= "000000000000000000000000";
		 i_in(6) <= "000000000000000000000000";
		 i_in(7) <= "000000000000000000000000";
		 i_in(8) <= "000000000000000000000000";
		 i_in(9) <= "000000000000000000000000";
		 i_in(10) <= "000000000000000000000000";
		 i_in(11) <= "000000000000000000000000";
		 i_in(12) <= "000000000000000000000000";
		 i_in(13) <= "000000000000000000000000";
		 i_in(14) <= "000000000000000000000000";
		 i_in(15) <= "000000000000000000000000";
	 
	 wait for 1*period;
	 TB_START <= '0';
	
	wait for 12*period;
	TB_START <= '1';
			
	 ---------------------- TEST 4 ---------------------- -1 -1 1 1 -1 -1 1 1 -1 -1 1 1 -1 -1 1 1 
		r_in(0) <= "100000000000000000000000";
		r_in(1) <= "100000000000000000000000";
		r_in(2) <= "011111111111111111111111";
		r_in(3) <= "011111111111111111111111";
		r_in(4) <= "100000000000000000000000";
		r_in(5) <= "100000000000000000000000";
		r_in(6) <= "011111111111111111111111";
		r_in(7) <= "011111111111111111111111";
		r_in(8) <= "100000000000000000000000";
		r_in(9) <= "100000000000000000000000";
		r_in(10) <= "011111111111111111111111";
		r_in(11) <= "011111111111111111111111";
		r_in(12) <= "100000000000000000000000";
		r_in(13) <= "100000000000000000000000";
		r_in(14) <= "011111111111111111111111";
		r_in(15) <= "011111111111111111111111";
		
		i_in(0) <= "000000000000000000000000";
		i_in(1) <= "000000000000000000000000";
		i_in(2) <= "000000000000000000000000";
		i_in(3) <= "000000000000000000000000";
		i_in(4) <= "000000000000000000000000";
		i_in(5) <= "000000000000000000000000";
		i_in(6) <= "000000000000000000000000";
		i_in(7) <= "000000000000000000000000";
		i_in(8) <= "000000000000000000000000";
		i_in(9) <= "000000000000000000000000";
		i_in(10) <= "000000000000000000000000";
		i_in(11) <= "000000000000000000000000";
		i_in(12) <= "000000000000000000000000";
		i_in(13) <= "000000000000000000000000";
		i_in(14) <= "000000000000000000000000";
		i_in(15) <= "000000000000000000000000";
	 
	 wait for 1*period;
	 TB_START <= '0';


	wait for 12*period;
	TB_START <= '1';
			
	 ---------------------- TEST 5 ---------------------- 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 -0.5 -0.5 -0.5 -0.5 -0.5 -0.5 -0.5
		r_in(0) <= "010000000000000000000000";
		r_in(1) <= "010000000000000000000000";
		r_in(2) <= "010000000000000000000000";
		r_in(3) <= "010000000000000000000000";
		r_in(4) <= "010000000000000000000000";
		r_in(5) <= "010000000000000000000000";
		r_in(6) <= "010000000000000000000000";
		r_in(7) <= "010000000000000000000000";
		r_in(8) <= "010000000000000000000000";
		r_in(9) <= "110000000000000000000000";
		r_in(10) <= "110000000000000000000000";
		r_in(11) <= "110000000000000000000000";
		r_in(12) <= "110000000000000000000000";
		r_in(13) <= "110000000000000000000000";
		r_in(14) <= "110000000000000000000000";
		r_in(15) <= "110000000000000000000000";
		
		i_in(0) <= "000000000000000000000000";
		i_in(1) <= "000000000000000000000000";
		i_in(2) <= "000000000000000000000000";
		i_in(3) <= "000000000000000000000000";
		i_in(4) <= "000000000000000000000000";
		i_in(5) <= "000000000000000000000000";
		i_in(6) <= "000000000000000000000000";
		i_in(7) <= "000000000000000000000000";
		i_in(8) <= "000000000000000000000000";
		i_in(9) <= "000000000000000000000000";
		i_in(10) <= "000000000000000000000000";
		i_in(11) <= "000000000000000000000000";
		i_in(12) <= "000000000000000000000000";
		i_in(13) <= "000000000000000000000000";
		i_in(14) <= "000000000000000000000000";
		i_in(15) <= "000000000000000000000000";
	 
	 wait for 1*period;
	 TB_START <= '0';

	wait for 12*period;
	TB_START <= '1';
			
	---------------------- TEST 6 ---------------------- 0 0 0 0 0 0 0 0 0.75 0 0 0 0 0 0 0
		r_in(0) <= "000000000000000000000000";
		r_in(1) <= "000000000000000000000000";
		r_in(2) <= "000000000000000000000000";
		r_in(3) <= "000000000000000000000000";
		r_in(4) <= "000000000000000000000000";
		r_in(5) <= "000000000000000000000000";
		r_in(6) <= "000000000000000000000000";
		r_in(7) <= "000000000000000000000000";
		r_in(8) <= "011000000000000000000000";
		r_in(9) <= "000000000000000000000000";
		r_in(10) <= "000000000000000000000000";
		r_in(11) <= "000000000000000000000000";
		r_in(12) <= "000000000000000000000000";
		r_in(13) <= "000000000000000000000000";
		r_in(14) <= "000000000000000000000000";
		r_in(15) <= "000000000000000000000000";
		
		i_in(0) <= "000000000000000000000000";
		i_in(1) <= "000000000000000000000000";
		i_in(2) <= "000000000000000000000000";
		i_in(3) <= "000000000000000000000000";
		i_in(4) <= "000000000000000000000000";
		i_in(5) <= "000000000000000000000000";
		i_in(6) <= "000000000000000000000000";
		i_in(7) <= "000000000000000000000000";
		i_in(8) <= "000000000000000000000000";
		i_in(9) <= "000000000000000000000000";
		i_in(10) <= "000000000000000000000000";
		i_in(11) <= "000000000000000000000000";
		i_in(12) <= "000000000000000000000000";
		i_in(13) <= "000000000000000000000000";
		i_in(14) <= "000000000000000000000000";
		i_in(15) <= "000000000000000000000000";
	 
	 wait for 1*period;
	 TB_START <= '0';
	 
	 wait for 12*period;
	TB_START <= '1';
			
	 ---------------------- TEST 7 ---------------------- 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5 0.5
		r_in(0) <= "010000000000000000000000";
		r_in(1) <= "010000000000000000000000";
		r_in(2) <= "010000000000000000000000";
		r_in(3) <= "010000000000000000000000";
		r_in(4) <= "010000000000000000000000";
		r_in(5) <= "010000000000000000000000";
		r_in(6) <= "010000000000000000000000";
		r_in(7) <= "010000000000000000000000";
		r_in(8) <= "010000000000000000000000";
		r_in(9) <= "010000000000000000000000";
		r_in(10) <= "010000000000000000000000";
		r_in(11) <= "010000000000000000000000";
		r_in(12) <= "010000000000000000000000";
		r_in(13) <= "010000000000000000000000";
		r_in(14) <= "010000000000000000000000";
		r_in(15) <= "010000000000000000000000";
		
		i_in(0) <= "000000000000000000000000";
		i_in(1) <= "000000000000000000000000";
		i_in(2) <= "000000000000000000000000";
		i_in(3) <= "000000000000000000000000";
		i_in(4) <= "000000000000000000000000";
		i_in(5) <= "000000000000000000000000";
		i_in(6) <= "000000000000000000000000";
		i_in(7) <= "000000000000000000000000";
		i_in(8) <= "000000000000000000000000";
		i_in(9) <= "000000000000000000000000";
		i_in(10) <= "000000000000000000000000";
		i_in(11) <= "000000000000000000000000";
		i_in(12) <= "000000000000000000000000";
		i_in(13) <= "000000000000000000000000";
		i_in(14) <= "000000000000000000000000";
		i_in(15) <= "000000000000000000000000";
	 
	 wait for 1*period;
	 TB_START <= '0';

	 wait;
        
    end process;

end behavioral;